LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;
entity sinelut_entity IS
	generic(
			lut_bit_width : integer := 8;
			data_width: integer := 16
	);
	port(
		phase_in      	: in unsigned(lut_bit_width-1 downto 0);
		a_clk      		: in std_logic;
		reset         	: in std_logic;
		data          	: out std_logic_vector(15 downto 0)
	);
end sinelut_entity;

architecture sinelut_entity_arch of sinelut_entity is 
--LUT
	type sine_lut is array (0 to (2**lut_bit_width)-1) of integer;
	constant sinedata:sine_lut:= (0,196,393,589,784,979,1174,1368,1561,1753,1944,2134,2322,2509,2695,2879,3061,3242,3420,3597,3771,3943,4113,4280,4445,4606,4766,4922,5075,5225,5372,5516,5657,5794,5928,6058,6184,6307,6426,6541,6652,6759,6862,6961,7055,7146,7232,7314,7391,7464,7532,7596,7656,7710,7760,7806,7846,7882,7913,7940,7961,7978,7990,7998,8000,7998,7990,7978,7961,7940,7913,7882,7846,7806,7760,7710,7656,7596,7532,7464,7391,7314,7232,7146,7055,6961,6862,6759,6652,6541,6426,6307,6184,6058,5928,5794,5657,5516,5372,5225,5075,4922,4766,4606,4445,4280,4113,3943,3771,3597,3420,3242,3061,2879,2695,2509,2322,2134,1944,1753,1561,1368,1174,979,784,589,393,196,0,-196,-393,-589,-784,-979,-1174,-1368,-1561,-1753,-1944,-2134,-2322,-2509,-2695,-2879,-3061,-3242,-3420,-3597,-3771,-3943,-4113,-4280,-4445,-4606,-4766,-4922,-5075,-5225,-5372,-5516,-5657,-5794,-5928,-6058,-6184,-6307,-6426,-6541,-6652,-6759,-6862,-6961,-7055,-7146,-7232,-7314,-7391,-7464,-7532,-7596,-7656,-7710,-7760,-7806,-7846,-7882,-7913,-7940,-7961,-7978,-7990,-7998,-8000,-7998,-7990,-7978,-7961,-7940,-7913,-7882,-7846,-7806,-7760,-7710,-7656,-7596,-7532,-7464,-7391,-7314,-7232,-7146,-7055,-6961,-6862,-6759,-6652,-6541,-6426,-6307,-6184,-6058,-5928,-5794,-5657,-5516,-5372,-5225,-5075,-4922,-4766,-4606,-4445,-4280,-4113,-3943,-3771,-3597,-3420,-3242,-3061,-2879,-2695,-2509,-2322,-2134,-1944,-1753,-1561,-1368,-1174,-979,-784,-589,-393,-196);
	signal 	sdata    : std_logic_vector(15 downto 0);
begin
	process(a_clk,reset)
		variable lutindex : integer range 0 to (2**lut_bit_width)-1 := 0;
	begin
		if reset = '0' then
			data <= (others => '0');
			lutindex := 0;
		elsif rising_edge(a_clk) then
			lutindex := to_integer(phase_in);
			sdata <= std_logic_vector(to_signed(sinedata(lutindex), data_width));
			data <= sdata;
		end if;	
	end process;
end architecture;