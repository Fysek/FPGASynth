LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;
entity trilut_entity IS
	generic(
			lut_bit_width : integer := 8;
			data_width: integer := 16
	);
	port(
		phase_in      	: in unsigned(lut_bit_width-1 downto 0);
		a_clk      		: in std_logic;
		reset         	: in std_logic;
		data          	: out std_logic_vector(15 downto 0)
	);
end trilut_entity;

architecture trilut_entity_arch of trilut_entity is 
--LUT
	type sine_lut is array (0 to (2**lut_bit_width)-1) of integer;
	constant sinedata:sine_lut:= (-7875,-7750,-7625,-7500,-7375,-7250,-7125,-7000,-6875,-6750,-6625,-6500,-6375,-6250,-6125,-6000,-5875,-5750,-5625,-5500,-5375,-5250,-5125,-5000,-4875,-4750,-4625,-4500,-4375,-4250,-4125,-4000,-3875,-3750,-3625,-3500,-3375,-3250,-3125,-3000,-2875,-2750,-2625,-2500,-2375,-2250,-2125,-2000,-1875,-1750,-1625,-1500,-1375,-1250,-1125,-1000,-875,-750,-625,-500,-375,-250,-125,0,125,250,375,500,625,750,875,1000,1125,1250,1375,1500,1625,1750,1875,2000,2125,2250,2375,2500,2625,2750,2875,3000,3125,3250,3375,3500,3625,3750,3875,4000,4125,4250,4375,4500,4625,4750,4875,5000,5125,5250,5375,5500,5625,5750,5875,6000,6125,6250,6375,6500,6625,6750,6875,7000,7125,7250,7375,7500,7625,7750,7875,8000,7875,7750,7625,7500,7375,7250,7125,7000,6875,6750,6625,6500,6375,6250,6125,6000,5875,5750,5625,5500,5375,5250,5125,5000,4875,4750,4625,4500,4375,4250,4125,4000,3875,3750,3625,3500,3375,3250,3125,3000,2875,2750,2625,2500,2375,2250,2125,2000,1875,1750,1625,1500,1375,1250,1125,1000,875,750,625,500,375,250,125,0,-125,-250,-375,-500,-625,-750,-875,-1000,-1125,-1250,-1375,-1500,-1625,-1750,-1875,-2000,-2125,-2250,-2375,-2500,-2625,-2750,-2875,-3000,-3125,-3250,-3375,-3500,-3625,-3750,-3875,-4000,-4125,-4250,-4375,-4500,-4625,-4750,-4875,-5000,-5125,-5250,-5375,-5500,-5625,-5750,-5875,-6000,-6125,-6250,-6375,-6500,-6625,-6750,-6875,-7000,-7125,-7250,-7375,-7500,-7625,-7750,-7875,-8000);
	signal 	sdata    : std_logic_vector(15 downto 0);
begin
	process(a_clk,reset)
		variable lutindex : integer range 0 to (2**lut_bit_width)-1 := 0;
	begin
		if reset = '0' then
			data <= (others => '0');
			lutindex := 0;
		elsif rising_edge(a_clk) then
			lutindex := to_integer(phase_in);
			sdata <= std_logic_vector(to_signed(sinedata(lutindex), data_width));
			data <= sdata; 
		end if;	
	end process;
end architecture;