LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;
ENTITY sawlut_entity IS
	generic(
			lut_bit_width : integer := 8;
			data_width: integer := 16
	);
	port(
		phase_in      : in unsigned(lut_bit_width-1 downto 0);
		a_clk      	: in std_logic;
		reset         : in std_logic;
		data          : out std_logic_vector(15 downto 0)
	);
end sawlut_entity;

architecture sawlut_entity_arch of sawlut_entity is 
--LUT
	type sine_lut is array (0 to (2**lut_bit_width)-1) of integer;
	constant sinedata:sine_lut:= (-7938,-7876,-7814,-7752,-7690,-7628,-7566,-7504,-7442,-7380,-7318,-7256,-7194,-7132,-7070,-7008,-6946,-6884,-6822,-6760,-6698,-6636,-6574,-6512,-6450,-6388,-6326,-6264,-6202,-6140,-6078,-6016,-5954,-5892,-5830,-5768,-5706,-5644,-5582,-5520,-5458,-5396,-5334,-5272,-5210,-5148,-5086,-5024,-4962,-4900,-4838,-4776,-4714,-4652,-4590,-4528,-4466,-4404,-4342,-4280,-4218,-4156,-4094,-4032,-3970,-3908,-3846,-3784,-3722,-3660,-3598,-3536,-3474,-3412,-3350,-3288,-3226,-3164,-3102,-3040,-2978,-2916,-2854,-2792,-2730,-2668,-2606,-2544,-2482,-2420,-2358,-2296,-2234,-2172,-2110,-2048,-1986,-1924,-1862,-1800,-1738,-1676,-1614,-1552,-1490,-1428,-1366,-1304,-1242,-1180,-1118,-1056,-994,-932,-870,-808,-746,-684,-622,-560,-498,-436,-374,-312,-250,-188,-126,-64,-2,60,122,184,246,308,370,432,494,556,618,680,742,804,866,928,990,1052,1114,1176,1238,1300,1362,1424,1486,1548,1610,1672,1734,1796,1858,1920,1982,2044,2106,2168,2230,2292,2354,2416,2478,2540,2602,2664,2726,2788,2850,2912,2974,3036,3098,3160,3222,3284,3346,3408,3470,3532,3594,3656,3718,3780,3842,3904,3966,4028,4090,4152,4214,4276,4338,4400,4462,4524,4586,4648,4710,4772,4834,4896,4958,5020,5082,5144,5206,5268,5330,5392,5454,5516,5578,5640,5702,5764,5826,5888,5950,6012,6074,6136,6198,6260,6322,6384,6446,6508,6570,6632,6694,6756,6818,6880,6942,7004,7066,7128,7190,7252,7314,7376,7438,7500,7562,7624,7686,7748,7810,7872);
	signal 	sdata    : std_logic_vector(15 downto 0);

begin
	process(a_clk,reset)
		variable lutindex : integer range 0 to (2**lut_bit_width)-1 := 0;
	begin
		if reset = '0' then
			data <= (others => '0');
			lutindex := 0;
		elsif rising_edge(a_clk) then
			lutindex := to_integer(phase_in);
			sdata <= std_logic_vector(to_signed(sinedata(lutindex), data_width));
			data <= sdata; 
		end if;	
	end process;
end architecture;