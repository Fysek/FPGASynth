module synthesizer (

	input logic clk,
	input logic uart_rx,
	output logic [2:0] datap,
	output logic [2:0] datan,
	output logic clkp,
	output logic clkn

)
;


endmodule